module tb_controller(output err);
  
	//inputs
	reg clk;
	reg rst_n;
	reg start;
        reg [2:0] opcode;
	reg [1:0] ALU_op;
 	reg [1:0] shift_op;
        reg Z;
	reg N;
	reg V;

	//outputs
        reg waiting;
        reg [1:0] reg_sel;
	reg [1:0] wb_sel;
	reg w_en;
       	reg en_A; 
	reg en_B;
	reg en_C;  
	reg en_status;
        reg sel_A;
	reg sel_B;

	reg error;
	assign err = error;

	parameter Rm = 2'b00;
	parameter Rd = 2'b01;
	parameter Rn = 2'b10;

	controller testBench(.clk, .rst_n, .start, .opcode, .ALU_op, .shift_op, .Z, .N, .V, .waiting, .reg_sel, .wb_sel, .w_en, .en_A, .en_B, .en_C, .en_status, .sel_A, .sel_B);



	initial begin
		forever begin
			clk = 1'b0;
			#10;
			clk = 1'b1;
			#10;
		end
	end



	initial begin
		error = 1'b0;
		//restart the fsm
		rst_n = 1'b0;
		
		#20;
		rst_n = 1'b1;


		//check move immediate
		start = 1'b1;
		opcode = 3'b110;
		ALU_op = 2'b10;
		
		#20;
		assert(w_en === 1'b1 && reg_sel === 2'b10 && wb_sel === 2'b10) $display("[PASS] MOV immediate");
     		else begin 
			$error("[FAIL] MOV immediate");
			error = 1;
		end


		
		//check move normal
		start = 1'b1;
		opcode = 3'b110;
		ALU_op = 2'b00;
		
		#20; //wait-> cycle 1 (1st)
		
		assert(reg_sel == Rm &&	en_A == 1'b0 && en_B == 1'b1) $display("[PASS] MOV normal cycle 1");
     		else begin 
			$error("[FAIL] MOV normal cycle 1");
			error = 1;
		end
		

		#20; //cycle 2 -> cycle 3

		assert(en_C == 1'b1 && sel_A == 1'b0 && sel_B == 1'b0) $display("[PASS] MOV normal cycle 3");
     		else begin 
			$error("[FAIL] MOV normal cycle 3");
			error = 1;
		end
		start = 1'b0;
		#20; //cycle 3 -> cycle 4

		assert(wb_sel == 2'b00 && w_en == 1'b1 && en_status == 1'b0) $display("[PASS] MOV normal cycle 4");
     		else begin 
			$error("[FAIL] MOV normal cycle 4");
			error = 1;
		end
	
		#20; //cycle 4 -> waiting state
		
		assert(waiting == 1'b1) $display("[PASS] MOV normal wait");
     		else begin 
			$error("[FAIL] MOV normal wait");
			error = 1;
		end


		//check ADD
		start = 1'b1;
		opcode = 3'b101;
		ALU_op = 2'b00;
		#20; 


		assert(reg_sel == Rn &&	en_A == 1'b1 && en_B == 1'b0) $display("[PASS] ADD cycle 1");
     		else begin 
			$error("[FAIL] ADD cycle 1");
			error = 1;
		end

		
		#20; //cycle 2

		assert(reg_sel == Rm &&	en_A == 1'b0 && en_B == 1'b1) $display("[PASS] ADD cycle 2");
     		else begin 
			$error("[FAIL] ADD cycle 2");
			error = 1;
		end

		start = 1'b0; //set start back to 0
		#20; //cycle 3
		
		assert(en_C == 1'b1 && sel_A == 1'b0 && sel_B == 1'b0 && en_status == 1'b1) $display("[PASS] ADD cycle 3");
     		else begin 
			$error("[FAIL] ADD cycle 3");
			error = 1;
		end
		
		#20; //cycle 4

		assert(wb_sel == 2'b00 && w_en == 1'b1 && en_status == 1'b0) $display("[PASS] ADD cycle 4");
     		else begin 
			$error("[FAIL] ADD cycle 4");
			error = 1;
		end


		#20; //wait state
		
		assert(waiting == 1'b1) $display("[PASS] ADD wait");
     		else begin 
			$error("[FAIL] ADD wait");
			error = 1;
		end

		//check CMP
		start = 1'b1;
		opcode = 3'b101;
		ALU_op = 2'b01;
		#20; 


		assert(reg_sel == Rn &&	en_A == 1'b1 && en_B == 1'b0) $display("[PASS] CMP cycle 1");
     		else begin 
			$error("[FAIL] CMP cycle 1");
			error = 1;
		end

		#20;

		assert(reg_sel == Rm &&	en_A == 1'b0 && en_B == 1'b1) $display("[PASS] CMP cycle 2");
     		else begin 
			$error("[FAIL] CMP cycle 2");
			error = 1;
		end

		start = 1'b0; //set start back to 0
		#20;

		assert(en_C == 1'b1 && sel_A == 1'b0 && sel_B == 1'b0 && en_status == 1'b1) $display("[PASS] CMP cycle 3");
     		else begin 
			$error("[FAIL] CMP cycle 3");
			error = 1;
		end
		
		#20;
		
		assert(waiting == 1'b1) $display("[PASS] CMP wait");
     		else begin 
			$error("[FAIL] CMP wait");
			error = 1;
		end
		
		//check AND
		start = 1'b1;
		opcode = 3'b101;
		ALU_op = 2'b10;
		#20; 

	
		assert(reg_sel == Rn &&	en_A == 1'b1 && en_B == 1'b0) $display("[PASS] AND cycle 1");
     		else begin 
			$error("[FAIL] AND cycle 1");
			error = 1;
		end

		#20; 

		assert(reg_sel == Rm &&	en_A == 1'b0 && en_B == 1'b1) $display("[PASS] AND cycle 2");
     		else begin 
			$error("[FAIL] AND cycle 2");
			error = 1;
		end

		start = 1'b0; //set start back to 0
		#20; //cycle 3
		
		assert(en_C == 1'b1 && sel_A == 1'b0 && sel_B == 1'b0 && en_status == 1'b1) $display("[PASS] AND cycle 3");
     		else begin 
			$error("[FAIL] AND cycle 3");
			error = 1;
		end
		
		#20; //cycle 4

		assert(wb_sel == 2'b00 && w_en == 1'b1 && en_status == 1'b0) $display("[PASS] AND cycle 4");
     		else begin 
			$error("[FAIL] AND cycle 4");
			error = 1;
		end


		#20; //wait state
		
		assert(waiting == 1'b1) $display("[PASS] AND wait");
     		else begin 
			$error("[FAIL] AND wait");
			error = 1;
		end


		//check mvn
		start = 1'b1;
		opcode = 3'b101;
		ALU_op = 2'b11;
		#20;

		assert(reg_sel == Rm &&	en_A == 1'b0 && en_B == 1'b1) $display("[PASS] MVN cycle 1");
     		else begin 
			$error("[FAIL] MVN cycle 1");
			error = 1;
		end

		#20;
		
		start = 1'b0;
		assert(en_C == 1'b1 && sel_A == 1'b0 && sel_B == 1'b0 && en_status == 1'b1) $display("[PASS] MVN cycle 3");
     		else begin 
			$error("[FAIL] MVN cycle 3");
			error = 1;
		end

		#20;

		assert(wb_sel == 2'b00 && w_en == 1'b1 && en_status == 1'b0) $display("[PASS] MVN cycle 4");
     		else begin 
			$error("[FAIL] MVN cycle 4");
			error = 1;
		end

		#20;
		
		assert(waiting == 1'b1) $display("[PASS] MVN wait");
     		else begin 
			$error("[FAIL] MVN wait");
			error = 1;
		end



	$stop;
	end
	
endmodule: tb_controller
